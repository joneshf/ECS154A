library verilog;
use verilog.vl_types.all;
entity project_01_vlg_check_tst is
    port(
        E               : in     vl_logic;
        N               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end project_01_vlg_check_tst;
