library verilog;
use verilog.vl_types.all;
entity EightBitAnd_vlg_check_tst is
    port(
        C               : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end EightBitAnd_vlg_check_tst;
