library verilog;
use verilog.vl_types.all;
entity OneBitFullAdder_vlg_vec_tst is
end OneBitFullAdder_vlg_vec_tst;
