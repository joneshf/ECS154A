library verilog;
use verilog.vl_types.all;
entity EightBitAnd_vlg_vec_tst is
end EightBitAnd_vlg_vec_tst;
