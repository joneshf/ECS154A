library verilog;
use verilog.vl_types.all;
entity EightBitNot_vlg_vec_tst is
end EightBitNot_vlg_vec_tst;
