library verilog;
use verilog.vl_types.all;
entity EightBitXor_vlg_vec_tst is
end EightBitXor_vlg_vec_tst;
