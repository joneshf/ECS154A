library verilog;
use verilog.vl_types.all;
entity compare_vlg_vec_tst is
end compare_vlg_vec_tst;
