library verilog;
use verilog.vl_types.all;
entity EightBitRot_vlg_vec_tst is
end EightBitRot_vlg_vec_tst;
