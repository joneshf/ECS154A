library verilog;
use verilog.vl_types.all;
entity gray_vlg_vec_tst is
end gray_vlg_vec_tst;
