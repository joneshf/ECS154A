library verilog;
use verilog.vl_types.all;
entity EightBitAdd_vlg_vec_tst is
end EightBitAdd_vlg_vec_tst;
