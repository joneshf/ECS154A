library verilog;
use verilog.vl_types.all;
entity FourBitcarryLookaheadAdder_vlg_vec_tst is
end FourBitcarryLookaheadAdder_vlg_vec_tst;
